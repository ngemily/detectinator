`ifndef _global_vh_
`define _global_vh_

`define DEBUG

`define MEM_SIZE 'h10_0000
`define WORD_SIZE 8
`define PIXEL_SIZE 24

`endif
