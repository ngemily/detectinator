`ifndef _global_vh_
`define _global_vh_

//`define DEBUG

`define MEM_SIZE 'h10_0000
`define C_TABLE_SIZE 255

`define WORD_SIZE 8
`define PIXEL_SIZE 24

`define IFILE "imgs/balloon.bmp"
`define OFILE "out/out.bmp"
`define CFILE "src/colors.txt"

`endif
