`ifndef _global_vh_
`define _global_vh_

//`define DEBUG

`define MEM_SIZE 'h10_0000
`define C_TABLE_SIZE 255

`define WORD_SIZE 8
`define MAX 255
`define MIN 0
`define PIXEL_SIZE 24

`define IFILE "imgs/alien.bmp"
`define OFILE "out/out.bmp"
`define CFILE "src/colors.txt"

`define FRAME_WIDTH 550     //0x226
`define FRAME_HEIGHT 303    // 0x12f

`define THRESHOLD 50

`endif
